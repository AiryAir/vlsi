`timescale 1ns / 1ps
module half_adder(
 input X,
 input Y,
 output C,
 output S
 );
xor x1(S,X,Y);
and n(C,X,Y);
 
endmodule
